-----------------------------------------------------------
--  Ver  :| Original Author   		:| Additional Author :| 
--  V1.0 :| Simon Doherty			   :| Eric Lunty        :| 
-----------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity sin_lut_effect is

port (
	clk      : in  std_logic;
	en       : in  std_logic;
	
	--Address inputs
	addr     : in  std_logic_vector(11 downto 0);
	
	--Sine outputs
	sin_out  : out std_logic_vector(11 downto 0));
end entity;


architecture rtl of sin_lut_effect is


type rom_type is array (0 to 4095) of std_logic_vector (11 downto 0);

constant SIN_ROM : rom_type :=

(
X"BFF",X"C01",X"C02",X"C04",X"C05",X"C07",X"C08",X"C0A",
X"C0C",X"C0D",X"C0F",X"C10",X"C12",X"C13",X"C15",X"C17",
X"C18",X"C1A",X"C1B",X"C1D",X"C1E",X"C20",X"C22",X"C23",
X"C25",X"C26",X"C28",X"C29",X"C2B",X"C2D",X"C2E",X"C30",
X"C31",X"C33",X"C34",X"C36",X"C38",X"C39",X"C3B",X"C3C",
X"C3E",X"C3F",X"C41",X"C42",X"C44",X"C46",X"C47",X"C49",
X"C4A",X"C4C",X"C4D",X"C4F",X"C51",X"C52",X"C54",X"C55",
X"C57",X"C58",X"C5A",X"C5C",X"C5D",X"C5F",X"C60",X"C62",
X"C63",X"C65",X"C66",X"C68",X"C6A",X"C6B",X"C6D",X"C6E",
X"C70",X"C71",X"C73",X"C75",X"C76",X"C78",X"C79",X"C7B",
X"C7C",X"C7E",X"C7F",X"C81",X"C83",X"C84",X"C86",X"C87",
X"C89",X"C8A",X"C8C",X"C8D",X"C8F",X"C91",X"C92",X"C94",
X"C95",X"C97",X"C98",X"C9A",X"C9B",X"C9D",X"C9F",X"CA0",
X"CA2",X"CA3",X"CA5",X"CA6",X"CA8",X"CA9",X"CAB",X"CAD",
X"CAE",X"CB0",X"CB1",X"CB3",X"CB4",X"CB6",X"CB7",X"CB9",
X"CBA",X"CBC",X"CBE",X"CBF",X"CC1",X"CC2",X"CC4",X"CC5",
X"CC7",X"CC8",X"CCA",X"CCB",X"CCD",X"CCE",X"CD0",X"CD2",
X"CD3",X"CD5",X"CD6",X"CD8",X"CD9",X"CDB",X"CDC",X"CDE",
X"CDF",X"CE1",X"CE2",X"CE4",X"CE5",X"CE7",X"CE9",X"CEA",
X"CEC",X"CED",X"CEF",X"CF0",X"CF2",X"CF3",X"CF5",X"CF6",
X"CF8",X"CF9",X"CFB",X"CFC",X"CFE",X"CFF",X"D01",X"D02",
X"D04",X"D06",X"D07",X"D09",X"D0A",X"D0C",X"D0D",X"D0F",
X"D10",X"D12",X"D13",X"D15",X"D16",X"D18",X"D19",X"D1B",
X"D1C",X"D1E",X"D1F",X"D21",X"D22",X"D24",X"D25",X"D27",
X"D28",X"D2A",X"D2B",X"D2D",X"D2E",X"D30",X"D31",X"D33",
X"D34",X"D36",X"D37",X"D39",X"D3A",X"D3C",X"D3D",X"D3F",
X"D40",X"D42",X"D43",X"D45",X"D46",X"D48",X"D49",X"D4B",
X"D4C",X"D4E",X"D4F",X"D51",X"D52",X"D54",X"D55",X"D56",
X"D58",X"D59",X"D5B",X"D5C",X"D5E",X"D5F",X"D61",X"D62",
X"D64",X"D65",X"D67",X"D68",X"D6A",X"D6B",X"D6D",X"D6E",
X"D70",X"D71",X"D72",X"D74",X"D75",X"D77",X"D78",X"D7A",
X"D7B",X"D7D",X"D7E",X"D80",X"D81",X"D83",X"D84",X"D85",
X"D87",X"D88",X"D8A",X"D8B",X"D8D",X"D8E",X"D90",X"D91",
X"D92",X"D94",X"D95",X"D97",X"D98",X"D9A",X"D9B",X"D9D",
X"D9E",X"D9F",X"DA1",X"DA2",X"DA4",X"DA5",X"DA7",X"DA8",
X"DA9",X"DAB",X"DAC",X"DAE",X"DAF",X"DB1",X"DB2",X"DB3",
X"DB5",X"DB6",X"DB8",X"DB9",X"DBA",X"DBC",X"DBD",X"DBF",
X"DC0",X"DC2",X"DC3",X"DC4",X"DC6",X"DC7",X"DC9",X"DCA",
X"DCB",X"DCD",X"DCE",X"DD0",X"DD1",X"DD2",X"DD4",X"DD5",
X"DD7",X"DD8",X"DD9",X"DDB",X"DDC",X"DDE",X"DDF",X"DE0",
X"DE2",X"DE3",X"DE4",X"DE6",X"DE7",X"DE9",X"DEA",X"DEB",
X"DED",X"DEE",X"DF0",X"DF1",X"DF2",X"DF4",X"DF5",X"DF6",
X"DF8",X"DF9",X"DFA",X"DFC",X"DFD",X"DFF",X"E00",X"E01",
X"E03",X"E04",X"E05",X"E07",X"E08",X"E09",X"E0B",X"E0C",
X"E0D",X"E0F",X"E10",X"E11",X"E13",X"E14",X"E16",X"E17",
X"E18",X"E1A",X"E1B",X"E1C",X"E1E",X"E1F",X"E20",X"E22",
X"E23",X"E24",X"E25",X"E27",X"E28",X"E29",X"E2B",X"E2C",
X"E2D",X"E2F",X"E30",X"E31",X"E33",X"E34",X"E35",X"E37",
X"E38",X"E39",X"E3B",X"E3C",X"E3D",X"E3E",X"E40",X"E41",
X"E42",X"E44",X"E45",X"E46",X"E47",X"E49",X"E4A",X"E4B",
X"E4D",X"E4E",X"E4F",X"E50",X"E52",X"E53",X"E54",X"E56",
X"E57",X"E58",X"E59",X"E5B",X"E5C",X"E5D",X"E5E",X"E60",
X"E61",X"E62",X"E64",X"E65",X"E66",X"E67",X"E69",X"E6A",
X"E6B",X"E6C",X"E6E",X"E6F",X"E70",X"E71",X"E73",X"E74",
X"E75",X"E76",X"E77",X"E79",X"E7A",X"E7B",X"E7C",X"E7E",
X"E7F",X"E80",X"E81",X"E83",X"E84",X"E85",X"E86",X"E87",
X"E89",X"E8A",X"E8B",X"E8C",X"E8D",X"E8F",X"E90",X"E91",
X"E92",X"E93",X"E95",X"E96",X"E97",X"E98",X"E99",X"E9B",
X"E9C",X"E9D",X"E9E",X"E9F",X"EA1",X"EA2",X"EA3",X"EA4",
X"EA5",X"EA6",X"EA8",X"EA9",X"EAA",X"EAB",X"EAC",X"EAE",
X"EAF",X"EB0",X"EB1",X"EB2",X"EB3",X"EB4",X"EB6",X"EB7",
X"EB8",X"EB9",X"EBA",X"EBB",X"EBD",X"EBE",X"EBF",X"EC0",
X"EC1",X"EC2",X"EC3",X"EC4",X"EC6",X"EC7",X"EC8",X"EC9",
X"ECA",X"ECB",X"ECC",X"ECE",X"ECF",X"ED0",X"ED1",X"ED2",
X"ED3",X"ED4",X"ED5",X"ED6",X"ED8",X"ED9",X"EDA",X"EDB",
X"EDC",X"EDD",X"EDE",X"EDF",X"EE0",X"EE1",X"EE2",X"EE4",
X"EE5",X"EE6",X"EE7",X"EE8",X"EE9",X"EEA",X"EEB",X"EEC",
X"EED",X"EEE",X"EEF",X"EF0",X"EF2",X"EF3",X"EF4",X"EF5",
X"EF6",X"EF7",X"EF8",X"EF9",X"EFA",X"EFB",X"EFC",X"EFD",
X"EFE",X"EFF",X"F00",X"F01",X"F02",X"F03",X"F04",X"F05",
X"F06",X"F07",X"F08",X"F09",X"F0A",X"F0B",X"F0D",X"F0E",
X"F0F",X"F10",X"F11",X"F12",X"F13",X"F14",X"F15",X"F16",
X"F17",X"F18",X"F19",X"F1A",X"F1B",X"F1C",X"F1D",X"F1D",
X"F1E",X"F1F",X"F20",X"F21",X"F22",X"F23",X"F24",X"F25",
X"F26",X"F27",X"F28",X"F29",X"F2A",X"F2B",X"F2C",X"F2D",
X"F2E",X"F2F",X"F30",X"F31",X"F32",X"F33",X"F34",X"F35",
X"F35",X"F36",X"F37",X"F38",X"F39",X"F3A",X"F3B",X"F3C",
X"F3D",X"F3E",X"F3F",X"F40",X"F41",X"F41",X"F42",X"F43",
X"F44",X"F45",X"F46",X"F47",X"F48",X"F49",X"F4A",X"F4A",
X"F4B",X"F4C",X"F4D",X"F4E",X"F4F",X"F50",X"F51",X"F52",
X"F52",X"F53",X"F54",X"F55",X"F56",X"F57",X"F58",X"F58",
X"F59",X"F5A",X"F5B",X"F5C",X"F5D",X"F5E",X"F5E",X"F5F",
X"F60",X"F61",X"F62",X"F63",X"F63",X"F64",X"F65",X"F66",
X"F67",X"F68",X"F68",X"F69",X"F6A",X"F6B",X"F6C",X"F6D",
X"F6D",X"F6E",X"F6F",X"F70",X"F71",X"F71",X"F72",X"F73",
X"F74",X"F74",X"F75",X"F76",X"F77",X"F78",X"F78",X"F79",
X"F7A",X"F7B",X"F7C",X"F7C",X"F7D",X"F7E",X"F7F",X"F7F",
X"F80",X"F81",X"F82",X"F82",X"F83",X"F84",X"F85",X"F85",
X"F86",X"F87",X"F88",X"F88",X"F89",X"F8A",X"F8A",X"F8B",
X"F8C",X"F8D",X"F8D",X"F8E",X"F8F",X"F90",X"F90",X"F91",
X"F92",X"F92",X"F93",X"F94",X"F94",X"F95",X"F96",X"F97",
X"F97",X"F98",X"F99",X"F99",X"F9A",X"F9B",X"F9B",X"F9C",
X"F9D",X"F9D",X"F9E",X"F9F",X"F9F",X"FA0",X"FA1",X"FA1",
X"FA2",X"FA3",X"FA3",X"FA4",X"FA5",X"FA5",X"FA6",X"FA7",
X"FA7",X"FA8",X"FA8",X"FA9",X"FAA",X"FAA",X"FAB",X"FAC",
X"FAC",X"FAD",X"FAD",X"FAE",X"FAF",X"FAF",X"FB0",X"FB0",
X"FB1",X"FB2",X"FB2",X"FB3",X"FB3",X"FB4",X"FB5",X"FB5",
X"FB6",X"FB6",X"FB7",X"FB8",X"FB8",X"FB9",X"FB9",X"FBA",
X"FBA",X"FBB",X"FBC",X"FBC",X"FBD",X"FBD",X"FBE",X"FBE",
X"FBF",X"FBF",X"FC0",X"FC0",X"FC1",X"FC2",X"FC2",X"FC3",
X"FC3",X"FC4",X"FC4",X"FC5",X"FC5",X"FC6",X"FC6",X"FC7",
X"FC7",X"FC8",X"FC8",X"FC9",X"FC9",X"FCA",X"FCA",X"FCB",
X"FCB",X"FCC",X"FCC",X"FCD",X"FCD",X"FCE",X"FCE",X"FCF",
X"FCF",X"FD0",X"FD0",X"FD1",X"FD1",X"FD2",X"FD2",X"FD2",
X"FD3",X"FD3",X"FD4",X"FD4",X"FD5",X"FD5",X"FD6",X"FD6",
X"FD6",X"FD7",X"FD7",X"FD8",X"FD8",X"FD9",X"FD9",X"FD9",
X"FDA",X"FDA",X"FDB",X"FDB",X"FDC",X"FDC",X"FDC",X"FDD",
X"FDD",X"FDE",X"FDE",X"FDE",X"FDF",X"FDF",X"FE0",X"FE0",
X"FE0",X"FE1",X"FE1",X"FE1",X"FE2",X"FE2",X"FE3",X"FE3",
X"FE3",X"FE4",X"FE4",X"FE4",X"FE5",X"FE5",X"FE5",X"FE6",
X"FE6",X"FE6",X"FE7",X"FE7",X"FE7",X"FE8",X"FE8",X"FE8",
X"FE9",X"FE9",X"FE9",X"FEA",X"FEA",X"FEA",X"FEB",X"FEB",
X"FEB",X"FEC",X"FEC",X"FEC",X"FED",X"FED",X"FED",X"FED",
X"FEE",X"FEE",X"FEE",X"FEF",X"FEF",X"FEF",X"FEF",X"FF0",
X"FF0",X"FF0",X"FF0",X"FF1",X"FF1",X"FF1",X"FF1",X"FF2",
X"FF2",X"FF2",X"FF2",X"FF3",X"FF3",X"FF3",X"FF3",X"FF4",
X"FF4",X"FF4",X"FF4",X"FF5",X"FF5",X"FF5",X"FF5",X"FF5",
X"FF6",X"FF6",X"FF6",X"FF6",X"FF7",X"FF7",X"FF7",X"FF7",
X"FF7",X"FF7",X"FF8",X"FF8",X"FF8",X"FF8",X"FF8",X"FF9",
X"FF9",X"FF9",X"FF9",X"FF9",X"FF9",X"FFA",X"FFA",X"FFA",
X"FFA",X"FFA",X"FFA",X"FFB",X"FFB",X"FFB",X"FFB",X"FFB",
X"FFB",X"FFB",X"FFB",X"FFC",X"FFC",X"FFC",X"FFC",X"FFC",
X"FFC",X"FFC",X"FFC",X"FFD",X"FFD",X"FFD",X"FFD",X"FFD",
X"FFD",X"FFD",X"FFD",X"FFD",X"FFD",X"FFE",X"FFE",X"FFE",
X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",
X"FFE",X"FFE",X"FFE",X"FFE",X"FFF",X"FFF",X"FFF",X"FFF",
X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",
X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",
X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",
X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",
X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFE",X"FFE",X"FFE",
X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",X"FFE",
X"FFE",X"FFE",X"FFE",X"FFE",X"FFD",X"FFD",X"FFD",X"FFD",
X"FFD",X"FFD",X"FFD",X"FFD",X"FFD",X"FFD",X"FFC",X"FFC",
X"FFC",X"FFC",X"FFC",X"FFC",X"FFC",X"FFC",X"FFB",X"FFB",
X"FFB",X"FFB",X"FFB",X"FFB",X"FFB",X"FFB",X"FFA",X"FFA",
X"FFA",X"FFA",X"FFA",X"FFA",X"FF9",X"FF9",X"FF9",X"FF9",
X"FF9",X"FF9",X"FF8",X"FF8",X"FF8",X"FF8",X"FF8",X"FF7",
X"FF7",X"FF7",X"FF7",X"FF7",X"FF7",X"FF6",X"FF6",X"FF6",
X"FF6",X"FF5",X"FF5",X"FF5",X"FF5",X"FF5",X"FF4",X"FF4",
X"FF4",X"FF4",X"FF3",X"FF3",X"FF3",X"FF3",X"FF2",X"FF2",
X"FF2",X"FF2",X"FF1",X"FF1",X"FF1",X"FF1",X"FF0",X"FF0",
X"FF0",X"FF0",X"FEF",X"FEF",X"FEF",X"FEF",X"FEE",X"FEE",
X"FEE",X"FED",X"FED",X"FED",X"FED",X"FEC",X"FEC",X"FEC",
X"FEB",X"FEB",X"FEB",X"FEA",X"FEA",X"FEA",X"FE9",X"FE9",
X"FE9",X"FE8",X"FE8",X"FE8",X"FE7",X"FE7",X"FE7",X"FE6",
X"FE6",X"FE6",X"FE5",X"FE5",X"FE5",X"FE4",X"FE4",X"FE4",
X"FE3",X"FE3",X"FE3",X"FE2",X"FE2",X"FE1",X"FE1",X"FE1",
X"FE0",X"FE0",X"FE0",X"FDF",X"FDF",X"FDE",X"FDE",X"FDE",
X"FDD",X"FDD",X"FDC",X"FDC",X"FDC",X"FDB",X"FDB",X"FDA",
X"FDA",X"FD9",X"FD9",X"FD9",X"FD8",X"FD8",X"FD7",X"FD7",
X"FD6",X"FD6",X"FD6",X"FD5",X"FD5",X"FD4",X"FD4",X"FD3",
X"FD3",X"FD2",X"FD2",X"FD2",X"FD1",X"FD1",X"FD0",X"FD0",
X"FCF",X"FCF",X"FCE",X"FCE",X"FCD",X"FCD",X"FCC",X"FCC",
X"FCB",X"FCB",X"FCA",X"FCA",X"FC9",X"FC9",X"FC8",X"FC8",
X"FC7",X"FC7",X"FC6",X"FC6",X"FC5",X"FC5",X"FC4",X"FC4",
X"FC3",X"FC3",X"FC2",X"FC2",X"FC1",X"FC0",X"FC0",X"FBF",
X"FBF",X"FBE",X"FBE",X"FBD",X"FBD",X"FBC",X"FBC",X"FBB",
X"FBA",X"FBA",X"FB9",X"FB9",X"FB8",X"FB8",X"FB7",X"FB6",
X"FB6",X"FB5",X"FB5",X"FB4",X"FB3",X"FB3",X"FB2",X"FB2",
X"FB1",X"FB0",X"FB0",X"FAF",X"FAF",X"FAE",X"FAD",X"FAD",
X"FAC",X"FAC",X"FAB",X"FAA",X"FAA",X"FA9",X"FA8",X"FA8",
X"FA7",X"FA7",X"FA6",X"FA5",X"FA5",X"FA4",X"FA3",X"FA3",
X"FA2",X"FA1",X"FA1",X"FA0",X"F9F",X"F9F",X"F9E",X"F9D",
X"F9D",X"F9C",X"F9B",X"F9B",X"F9A",X"F99",X"F99",X"F98",
X"F97",X"F97",X"F96",X"F95",X"F94",X"F94",X"F93",X"F92",
X"F92",X"F91",X"F90",X"F90",X"F8F",X"F8E",X"F8D",X"F8D",
X"F8C",X"F8B",X"F8A",X"F8A",X"F89",X"F88",X"F88",X"F87",
X"F86",X"F85",X"F85",X"F84",X"F83",X"F82",X"F82",X"F81",
X"F80",X"F7F",X"F7F",X"F7E",X"F7D",X"F7C",X"F7C",X"F7B",
X"F7A",X"F79",X"F78",X"F78",X"F77",X"F76",X"F75",X"F74",
X"F74",X"F73",X"F72",X"F71",X"F71",X"F70",X"F6F",X"F6E",
X"F6D",X"F6D",X"F6C",X"F6B",X"F6A",X"F69",X"F68",X"F68",
X"F67",X"F66",X"F65",X"F64",X"F63",X"F63",X"F62",X"F61",
X"F60",X"F5F",X"F5E",X"F5E",X"F5D",X"F5C",X"F5B",X"F5A",
X"F59",X"F58",X"F58",X"F57",X"F56",X"F55",X"F54",X"F53",
X"F52",X"F52",X"F51",X"F50",X"F4F",X"F4E",X"F4D",X"F4C",
X"F4B",X"F4A",X"F4A",X"F49",X"F48",X"F47",X"F46",X"F45",
X"F44",X"F43",X"F42",X"F41",X"F41",X"F40",X"F3F",X"F3E",
X"F3D",X"F3C",X"F3B",X"F3A",X"F39",X"F38",X"F37",X"F36",
X"F35",X"F35",X"F34",X"F33",X"F32",X"F31",X"F30",X"F2F",
X"F2E",X"F2D",X"F2C",X"F2B",X"F2A",X"F29",X"F28",X"F27",
X"F26",X"F25",X"F24",X"F23",X"F22",X"F21",X"F20",X"F1F",
X"F1E",X"F1D",X"F1D",X"F1C",X"F1B",X"F1A",X"F19",X"F18",
X"F17",X"F16",X"F15",X"F14",X"F13",X"F12",X"F11",X"F10",
X"F0F",X"F0E",X"F0D",X"F0B",X"F0A",X"F09",X"F08",X"F07",
X"F06",X"F05",X"F04",X"F03",X"F02",X"F01",X"F00",X"EFF",
X"EFE",X"EFD",X"EFC",X"EFB",X"EFA",X"EF9",X"EF8",X"EF7",
X"EF6",X"EF5",X"EF4",X"EF3",X"EF2",X"EF0",X"EEF",X"EEE",
X"EED",X"EEC",X"EEB",X"EEA",X"EE9",X"EE8",X"EE7",X"EE6",
X"EE5",X"EE4",X"EE2",X"EE1",X"EE0",X"EDF",X"EDE",X"EDD",
X"EDC",X"EDB",X"EDA",X"ED9",X"ED8",X"ED6",X"ED5",X"ED4",
X"ED3",X"ED2",X"ED1",X"ED0",X"ECF",X"ECE",X"ECC",X"ECB",
X"ECA",X"EC9",X"EC8",X"EC7",X"EC6",X"EC4",X"EC3",X"EC2",
X"EC1",X"EC0",X"EBF",X"EBE",X"EBD",X"EBB",X"EBA",X"EB9",
X"EB8",X"EB7",X"EB6",X"EB4",X"EB3",X"EB2",X"EB1",X"EB0",
X"EAF",X"EAE",X"EAC",X"EAB",X"EAA",X"EA9",X"EA8",X"EA6",
X"EA5",X"EA4",X"EA3",X"EA2",X"EA1",X"E9F",X"E9E",X"E9D",
X"E9C",X"E9B",X"E99",X"E98",X"E97",X"E96",X"E95",X"E93",
X"E92",X"E91",X"E90",X"E8F",X"E8D",X"E8C",X"E8B",X"E8A",
X"E89",X"E87",X"E86",X"E85",X"E84",X"E83",X"E81",X"E80",
X"E7F",X"E7E",X"E7C",X"E7B",X"E7A",X"E79",X"E77",X"E76",
X"E75",X"E74",X"E73",X"E71",X"E70",X"E6F",X"E6E",X"E6C",
X"E6B",X"E6A",X"E69",X"E67",X"E66",X"E65",X"E64",X"E62",
X"E61",X"E60",X"E5E",X"E5D",X"E5C",X"E5B",X"E59",X"E58",
X"E57",X"E56",X"E54",X"E53",X"E52",X"E50",X"E4F",X"E4E",
X"E4D",X"E4B",X"E4A",X"E49",X"E47",X"E46",X"E45",X"E44",
X"E42",X"E41",X"E40",X"E3E",X"E3D",X"E3C",X"E3B",X"E39",
X"E38",X"E37",X"E35",X"E34",X"E33",X"E31",X"E30",X"E2F",
X"E2D",X"E2C",X"E2B",X"E29",X"E28",X"E27",X"E25",X"E24",
X"E23",X"E22",X"E20",X"E1F",X"E1E",X"E1C",X"E1B",X"E1A",
X"E18",X"E17",X"E16",X"E14",X"E13",X"E11",X"E10",X"E0F",
X"E0D",X"E0C",X"E0B",X"E09",X"E08",X"E07",X"E05",X"E04",
X"E03",X"E01",X"E00",X"DFF",X"DFD",X"DFC",X"DFA",X"DF9",
X"DF8",X"DF6",X"DF5",X"DF4",X"DF2",X"DF1",X"DF0",X"DEE",
X"DED",X"DEB",X"DEA",X"DE9",X"DE7",X"DE6",X"DE4",X"DE3",
X"DE2",X"DE0",X"DDF",X"DDE",X"DDC",X"DDB",X"DD9",X"DD8",
X"DD7",X"DD5",X"DD4",X"DD2",X"DD1",X"DD0",X"DCE",X"DCD",
X"DCB",X"DCA",X"DC9",X"DC7",X"DC6",X"DC4",X"DC3",X"DC2",
X"DC0",X"DBF",X"DBD",X"DBC",X"DBA",X"DB9",X"DB8",X"DB6",
X"DB5",X"DB3",X"DB2",X"DB1",X"DAF",X"DAE",X"DAC",X"DAB",
X"DA9",X"DA8",X"DA7",X"DA5",X"DA4",X"DA2",X"DA1",X"D9F",
X"D9E",X"D9D",X"D9B",X"D9A",X"D98",X"D97",X"D95",X"D94",
X"D92",X"D91",X"D90",X"D8E",X"D8D",X"D8B",X"D8A",X"D88",
X"D87",X"D85",X"D84",X"D83",X"D81",X"D80",X"D7E",X"D7D",
X"D7B",X"D7A",X"D78",X"D77",X"D75",X"D74",X"D72",X"D71",
X"D70",X"D6E",X"D6D",X"D6B",X"D6A",X"D68",X"D67",X"D65",
X"D64",X"D62",X"D61",X"D5F",X"D5E",X"D5C",X"D5B",X"D59",
X"D58",X"D56",X"D55",X"D54",X"D52",X"D51",X"D4F",X"D4E",
X"D4C",X"D4B",X"D49",X"D48",X"D46",X"D45",X"D43",X"D42",
X"D40",X"D3F",X"D3D",X"D3C",X"D3A",X"D39",X"D37",X"D36",
X"D34",X"D33",X"D31",X"D30",X"D2E",X"D2D",X"D2B",X"D2A",
X"D28",X"D27",X"D25",X"D24",X"D22",X"D21",X"D1F",X"D1E",
X"D1C",X"D1B",X"D19",X"D18",X"D16",X"D15",X"D13",X"D12",
X"D10",X"D0F",X"D0D",X"D0C",X"D0A",X"D09",X"D07",X"D06",
X"D04",X"D02",X"D01",X"CFF",X"CFE",X"CFC",X"CFB",X"CF9",
X"CF8",X"CF6",X"CF5",X"CF3",X"CF2",X"CF0",X"CEF",X"CED",
X"CEC",X"CEA",X"CE9",X"CE7",X"CE5",X"CE4",X"CE2",X"CE1",
X"CDF",X"CDE",X"CDC",X"CDB",X"CD9",X"CD8",X"CD6",X"CD5",
X"CD3",X"CD2",X"CD0",X"CCE",X"CCD",X"CCB",X"CCA",X"CC8",
X"CC7",X"CC5",X"CC4",X"CC2",X"CC1",X"CBF",X"CBE",X"CBC",
X"CBA",X"CB9",X"CB7",X"CB6",X"CB4",X"CB3",X"CB1",X"CB0",
X"CAE",X"CAD",X"CAB",X"CA9",X"CA8",X"CA6",X"CA5",X"CA3",
X"CA2",X"CA0",X"C9F",X"C9D",X"C9B",X"C9A",X"C98",X"C97",
X"C95",X"C94",X"C92",X"C91",X"C8F",X"C8D",X"C8C",X"C8A",
X"C89",X"C87",X"C86",X"C84",X"C83",X"C81",X"C7F",X"C7E",
X"C7C",X"C7B",X"C79",X"C78",X"C76",X"C75",X"C73",X"C71",
X"C70",X"C6E",X"C6D",X"C6B",X"C6A",X"C68",X"C66",X"C65",
X"C63",X"C62",X"C60",X"C5F",X"C5D",X"C5C",X"C5A",X"C58",
X"C57",X"C55",X"C54",X"C52",X"C51",X"C4F",X"C4D",X"C4C",
X"C4A",X"C49",X"C47",X"C46",X"C44",X"C42",X"C41",X"C3F",
X"C3E",X"C3C",X"C3B",X"C39",X"C38",X"C36",X"C34",X"C33",
X"C31",X"C30",X"C2E",X"C2D",X"C2B",X"C29",X"C28",X"C26",
X"C25",X"C23",X"C22",X"C20",X"C1E",X"C1D",X"C1B",X"C1A",
X"C18",X"C17",X"C15",X"C13",X"C12",X"C10",X"C0F",X"C0D",
X"C0C",X"C0A",X"C08",X"C07",X"C05",X"C04",X"C02",X"C01",
X"BFF",X"BFD",X"BFC",X"BFA",X"BF9",X"BF7",X"BF6",X"BF4",
X"BF2",X"BF1",X"BEF",X"BEE",X"BEC",X"BEB",X"BE9",X"BE7",
X"BE6",X"BE4",X"BE3",X"BE1",X"BE0",X"BDE",X"BDC",X"BDB",
X"BD9",X"BD8",X"BD6",X"BD5",X"BD3",X"BD1",X"BD0",X"BCE",
X"BCD",X"BCB",X"BCA",X"BC8",X"BC6",X"BC5",X"BC3",X"BC2",
X"BC0",X"BBF",X"BBD",X"BBC",X"BBA",X"BB8",X"BB7",X"BB5",
X"BB4",X"BB2",X"BB1",X"BAF",X"BAD",X"BAC",X"BAA",X"BA9",
X"BA7",X"BA6",X"BA4",X"BA2",X"BA1",X"B9F",X"B9E",X"B9C",
X"B9B",X"B99",X"B98",X"B96",X"B94",X"B93",X"B91",X"B90",
X"B8E",X"B8D",X"B8B",X"B89",X"B88",X"B86",X"B85",X"B83",
X"B82",X"B80",X"B7F",X"B7D",X"B7B",X"B7A",X"B78",X"B77",
X"B75",X"B74",X"B72",X"B71",X"B6F",X"B6D",X"B6C",X"B6A",
X"B69",X"B67",X"B66",X"B64",X"B63",X"B61",X"B5F",X"B5E",
X"B5C",X"B5B",X"B59",X"B58",X"B56",X"B55",X"B53",X"B51",
X"B50",X"B4E",X"B4D",X"B4B",X"B4A",X"B48",X"B47",X"B45",
X"B44",X"B42",X"B40",X"B3F",X"B3D",X"B3C",X"B3A",X"B39",
X"B37",X"B36",X"B34",X"B33",X"B31",X"B30",X"B2E",X"B2C",
X"B2B",X"B29",X"B28",X"B26",X"B25",X"B23",X"B22",X"B20",
X"B1F",X"B1D",X"B1C",X"B1A",X"B19",X"B17",X"B15",X"B14",
X"B12",X"B11",X"B0F",X"B0E",X"B0C",X"B0B",X"B09",X"B08",
X"B06",X"B05",X"B03",X"B02",X"B00",X"AFF",X"AFD",X"AFC",
X"AFA",X"AF8",X"AF7",X"AF5",X"AF4",X"AF2",X"AF1",X"AEF",
X"AEE",X"AEC",X"AEB",X"AE9",X"AE8",X"AE6",X"AE5",X"AE3",
X"AE2",X"AE0",X"ADF",X"ADD",X"ADC",X"ADA",X"AD9",X"AD7",
X"AD6",X"AD4",X"AD3",X"AD1",X"AD0",X"ACE",X"ACD",X"ACB",
X"ACA",X"AC8",X"AC7",X"AC5",X"AC4",X"AC2",X"AC1",X"ABF",
X"ABE",X"ABC",X"ABB",X"AB9",X"AB8",X"AB6",X"AB5",X"AB3",
X"AB2",X"AB0",X"AAF",X"AAD",X"AAC",X"AAA",X"AA9",X"AA8",
X"AA6",X"AA5",X"AA3",X"AA2",X"AA0",X"A9F",X"A9D",X"A9C",
X"A9A",X"A99",X"A97",X"A96",X"A94",X"A93",X"A91",X"A90",
X"A8E",X"A8D",X"A8C",X"A8A",X"A89",X"A87",X"A86",X"A84",
X"A83",X"A81",X"A80",X"A7E",X"A7D",X"A7B",X"A7A",X"A79",
X"A77",X"A76",X"A74",X"A73",X"A71",X"A70",X"A6E",X"A6D",
X"A6C",X"A6A",X"A69",X"A67",X"A66",X"A64",X"A63",X"A61",
X"A60",X"A5F",X"A5D",X"A5C",X"A5A",X"A59",X"A57",X"A56",
X"A55",X"A53",X"A52",X"A50",X"A4F",X"A4D",X"A4C",X"A4B",
X"A49",X"A48",X"A46",X"A45",X"A44",X"A42",X"A41",X"A3F",
X"A3E",X"A3C",X"A3B",X"A3A",X"A38",X"A37",X"A35",X"A34",
X"A33",X"A31",X"A30",X"A2E",X"A2D",X"A2C",X"A2A",X"A29",
X"A27",X"A26",X"A25",X"A23",X"A22",X"A20",X"A1F",X"A1E",
X"A1C",X"A1B",X"A1A",X"A18",X"A17",X"A15",X"A14",X"A13",
X"A11",X"A10",X"A0E",X"A0D",X"A0C",X"A0A",X"A09",X"A08",
X"A06",X"A05",X"A04",X"A02",X"A01",X"9FF",X"9FE",X"9FD",
X"9FB",X"9FA",X"9F9",X"9F7",X"9F6",X"9F5",X"9F3",X"9F2",
X"9F1",X"9EF",X"9EE",X"9ED",X"9EB",X"9EA",X"9E8",X"9E7",
X"9E6",X"9E4",X"9E3",X"9E2",X"9E0",X"9DF",X"9DE",X"9DC",
X"9DB",X"9DA",X"9D9",X"9D7",X"9D6",X"9D5",X"9D3",X"9D2",
X"9D1",X"9CF",X"9CE",X"9CD",X"9CB",X"9CA",X"9C9",X"9C7",
X"9C6",X"9C5",X"9C3",X"9C2",X"9C1",X"9C0",X"9BE",X"9BD",
X"9BC",X"9BA",X"9B9",X"9B8",X"9B7",X"9B5",X"9B4",X"9B3",
X"9B1",X"9B0",X"9AF",X"9AE",X"9AC",X"9AB",X"9AA",X"9A8",
X"9A7",X"9A6",X"9A5",X"9A3",X"9A2",X"9A1",X"9A0",X"99E",
X"99D",X"99C",X"99A",X"999",X"998",X"997",X"995",X"994",
X"993",X"992",X"990",X"98F",X"98E",X"98D",X"98B",X"98A",
X"989",X"988",X"987",X"985",X"984",X"983",X"982",X"980",
X"97F",X"97E",X"97D",X"97B",X"97A",X"979",X"978",X"977",
X"975",X"974",X"973",X"972",X"971",X"96F",X"96E",X"96D",
X"96C",X"96B",X"969",X"968",X"967",X"966",X"965",X"963",
X"962",X"961",X"960",X"95F",X"95D",X"95C",X"95B",X"95A",
X"959",X"958",X"956",X"955",X"954",X"953",X"952",X"950",
X"94F",X"94E",X"94D",X"94C",X"94B",X"94A",X"948",X"947",
X"946",X"945",X"944",X"943",X"941",X"940",X"93F",X"93E",
X"93D",X"93C",X"93B",X"93A",X"938",X"937",X"936",X"935",
X"934",X"933",X"932",X"930",X"92F",X"92E",X"92D",X"92C",
X"92B",X"92A",X"929",X"928",X"926",X"925",X"924",X"923",
X"922",X"921",X"920",X"91F",X"91E",X"91D",X"91C",X"91A",
X"919",X"918",X"917",X"916",X"915",X"914",X"913",X"912",
X"911",X"910",X"90F",X"90E",X"90C",X"90B",X"90A",X"909",
X"908",X"907",X"906",X"905",X"904",X"903",X"902",X"901",
X"900",X"8FF",X"8FE",X"8FD",X"8FC",X"8FB",X"8FA",X"8F9",
X"8F8",X"8F7",X"8F6",X"8F5",X"8F4",X"8F3",X"8F1",X"8F0",
X"8EF",X"8EE",X"8ED",X"8EC",X"8EB",X"8EA",X"8E9",X"8E8",
X"8E7",X"8E6",X"8E5",X"8E4",X"8E3",X"8E2",X"8E1",X"8E1",
X"8E0",X"8DF",X"8DE",X"8DD",X"8DC",X"8DB",X"8DA",X"8D9",
X"8D8",X"8D7",X"8D6",X"8D5",X"8D4",X"8D3",X"8D2",X"8D1",
X"8D0",X"8CF",X"8CE",X"8CD",X"8CC",X"8CB",X"8CA",X"8C9",
X"8C9",X"8C8",X"8C7",X"8C6",X"8C5",X"8C4",X"8C3",X"8C2",
X"8C1",X"8C0",X"8BF",X"8BE",X"8BD",X"8BD",X"8BC",X"8BB",
X"8BA",X"8B9",X"8B8",X"8B7",X"8B6",X"8B5",X"8B4",X"8B4",
X"8B3",X"8B2",X"8B1",X"8B0",X"8AF",X"8AE",X"8AD",X"8AC",
X"8AC",X"8AB",X"8AA",X"8A9",X"8A8",X"8A7",X"8A6",X"8A6",
X"8A5",X"8A4",X"8A3",X"8A2",X"8A1",X"8A0",X"8A0",X"89F",
X"89E",X"89D",X"89C",X"89B",X"89B",X"89A",X"899",X"898",
X"897",X"896",X"896",X"895",X"894",X"893",X"892",X"891",
X"891",X"890",X"88F",X"88E",X"88D",X"88D",X"88C",X"88B",
X"88A",X"88A",X"889",X"888",X"887",X"886",X"886",X"885",
X"884",X"883",X"882",X"882",X"881",X"880",X"87F",X"87F",
X"87E",X"87D",X"87C",X"87C",X"87B",X"87A",X"879",X"879",
X"878",X"877",X"876",X"876",X"875",X"874",X"874",X"873",
X"872",X"871",X"871",X"870",X"86F",X"86E",X"86E",X"86D",
X"86C",X"86C",X"86B",X"86A",X"86A",X"869",X"868",X"867",
X"867",X"866",X"865",X"865",X"864",X"863",X"863",X"862",
X"861",X"861",X"860",X"85F",X"85F",X"85E",X"85D",X"85D",
X"85C",X"85B",X"85B",X"85A",X"859",X"859",X"858",X"857",
X"857",X"856",X"856",X"855",X"854",X"854",X"853",X"852",
X"852",X"851",X"851",X"850",X"84F",X"84F",X"84E",X"84E",
X"84D",X"84C",X"84C",X"84B",X"84B",X"84A",X"849",X"849",
X"848",X"848",X"847",X"846",X"846",X"845",X"845",X"844",
X"844",X"843",X"842",X"842",X"841",X"841",X"840",X"840",
X"83F",X"83F",X"83E",X"83E",X"83D",X"83C",X"83C",X"83B",
X"83B",X"83A",X"83A",X"839",X"839",X"838",X"838",X"837",
X"837",X"836",X"836",X"835",X"835",X"834",X"834",X"833",
X"833",X"832",X"832",X"831",X"831",X"830",X"830",X"82F",
X"82F",X"82E",X"82E",X"82D",X"82D",X"82C",X"82C",X"82C",
X"82B",X"82B",X"82A",X"82A",X"829",X"829",X"828",X"828",
X"828",X"827",X"827",X"826",X"826",X"825",X"825",X"825",
X"824",X"824",X"823",X"823",X"822",X"822",X"822",X"821",
X"821",X"820",X"820",X"820",X"81F",X"81F",X"81E",X"81E",
X"81E",X"81D",X"81D",X"81D",X"81C",X"81C",X"81B",X"81B",
X"81B",X"81A",X"81A",X"81A",X"819",X"819",X"819",X"818",
X"818",X"818",X"817",X"817",X"817",X"816",X"816",X"816",
X"815",X"815",X"815",X"814",X"814",X"814",X"813",X"813",
X"813",X"812",X"812",X"812",X"811",X"811",X"811",X"811",
X"810",X"810",X"810",X"80F",X"80F",X"80F",X"80F",X"80E",
X"80E",X"80E",X"80E",X"80D",X"80D",X"80D",X"80D",X"80C",
X"80C",X"80C",X"80C",X"80B",X"80B",X"80B",X"80B",X"80A",
X"80A",X"80A",X"80A",X"809",X"809",X"809",X"809",X"809",
X"808",X"808",X"808",X"808",X"807",X"807",X"807",X"807",
X"807",X"807",X"806",X"806",X"806",X"806",X"806",X"805",
X"805",X"805",X"805",X"805",X"805",X"804",X"804",X"804",
X"804",X"804",X"804",X"803",X"803",X"803",X"803",X"803",
X"803",X"803",X"803",X"802",X"802",X"802",X"802",X"802",
X"802",X"802",X"802",X"801",X"801",X"801",X"801",X"801",
X"801",X"801",X"801",X"801",X"801",X"800",X"800",X"800",
X"800",X"800",X"800",X"800",X"800",X"800",X"800",X"800",
X"800",X"800",X"800",X"800",X"7FF",X"7FF",X"7FF",X"7FF",
X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",
X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",
X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",
X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",
X"7FF",X"7FF",X"7FF",X"7FF",X"7FF",X"800",X"800",X"800",
X"800",X"800",X"800",X"800",X"800",X"800",X"800",X"800",
X"800",X"800",X"800",X"800",X"801",X"801",X"801",X"801",
X"801",X"801",X"801",X"801",X"801",X"801",X"802",X"802",
X"802",X"802",X"802",X"802",X"802",X"802",X"803",X"803",
X"803",X"803",X"803",X"803",X"803",X"803",X"804",X"804",
X"804",X"804",X"804",X"804",X"805",X"805",X"805",X"805",
X"805",X"805",X"806",X"806",X"806",X"806",X"806",X"807",
X"807",X"807",X"807",X"807",X"807",X"808",X"808",X"808",
X"808",X"809",X"809",X"809",X"809",X"809",X"80A",X"80A",
X"80A",X"80A",X"80B",X"80B",X"80B",X"80B",X"80C",X"80C",
X"80C",X"80C",X"80D",X"80D",X"80D",X"80D",X"80E",X"80E",
X"80E",X"80E",X"80F",X"80F",X"80F",X"80F",X"810",X"810",
X"810",X"811",X"811",X"811",X"811",X"812",X"812",X"812",
X"813",X"813",X"813",X"814",X"814",X"814",X"815",X"815",
X"815",X"816",X"816",X"816",X"817",X"817",X"817",X"818",
X"818",X"818",X"819",X"819",X"819",X"81A",X"81A",X"81A",
X"81B",X"81B",X"81B",X"81C",X"81C",X"81D",X"81D",X"81D",
X"81E",X"81E",X"81E",X"81F",X"81F",X"820",X"820",X"820",
X"821",X"821",X"822",X"822",X"822",X"823",X"823",X"824",
X"824",X"825",X"825",X"825",X"826",X"826",X"827",X"827",
X"828",X"828",X"828",X"829",X"829",X"82A",X"82A",X"82B",
X"82B",X"82C",X"82C",X"82C",X"82D",X"82D",X"82E",X"82E",
X"82F",X"82F",X"830",X"830",X"831",X"831",X"832",X"832",
X"833",X"833",X"834",X"834",X"835",X"835",X"836",X"836",
X"837",X"837",X"838",X"838",X"839",X"839",X"83A",X"83A",
X"83B",X"83B",X"83C",X"83C",X"83D",X"83E",X"83E",X"83F",
X"83F",X"840",X"840",X"841",X"841",X"842",X"842",X"843",
X"844",X"844",X"845",X"845",X"846",X"846",X"847",X"848",
X"848",X"849",X"849",X"84A",X"84B",X"84B",X"84C",X"84C",
X"84D",X"84E",X"84E",X"84F",X"84F",X"850",X"851",X"851",
X"852",X"852",X"853",X"854",X"854",X"855",X"856",X"856",
X"857",X"857",X"858",X"859",X"859",X"85A",X"85B",X"85B",
X"85C",X"85D",X"85D",X"85E",X"85F",X"85F",X"860",X"861",
X"861",X"862",X"863",X"863",X"864",X"865",X"865",X"866",
X"867",X"867",X"868",X"869",X"86A",X"86A",X"86B",X"86C",
X"86C",X"86D",X"86E",X"86E",X"86F",X"870",X"871",X"871",
X"872",X"873",X"874",X"874",X"875",X"876",X"876",X"877",
X"878",X"879",X"879",X"87A",X"87B",X"87C",X"87C",X"87D",
X"87E",X"87F",X"87F",X"880",X"881",X"882",X"882",X"883",
X"884",X"885",X"886",X"886",X"887",X"888",X"889",X"88A",
X"88A",X"88B",X"88C",X"88D",X"88D",X"88E",X"88F",X"890",
X"891",X"891",X"892",X"893",X"894",X"895",X"896",X"896",
X"897",X"898",X"899",X"89A",X"89B",X"89B",X"89C",X"89D",
X"89E",X"89F",X"8A0",X"8A0",X"8A1",X"8A2",X"8A3",X"8A4",
X"8A5",X"8A6",X"8A6",X"8A7",X"8A8",X"8A9",X"8AA",X"8AB",
X"8AC",X"8AC",X"8AD",X"8AE",X"8AF",X"8B0",X"8B1",X"8B2",
X"8B3",X"8B4",X"8B4",X"8B5",X"8B6",X"8B7",X"8B8",X"8B9",
X"8BA",X"8BB",X"8BC",X"8BD",X"8BD",X"8BE",X"8BF",X"8C0",
X"8C1",X"8C2",X"8C3",X"8C4",X"8C5",X"8C6",X"8C7",X"8C8",
X"8C9",X"8C9",X"8CA",X"8CB",X"8CC",X"8CD",X"8CE",X"8CF",
X"8D0",X"8D1",X"8D2",X"8D3",X"8D4",X"8D5",X"8D6",X"8D7",
X"8D8",X"8D9",X"8DA",X"8DB",X"8DC",X"8DD",X"8DE",X"8DF",
X"8E0",X"8E1",X"8E1",X"8E2",X"8E3",X"8E4",X"8E5",X"8E6",
X"8E7",X"8E8",X"8E9",X"8EA",X"8EB",X"8EC",X"8ED",X"8EE",
X"8EF",X"8F0",X"8F1",X"8F3",X"8F4",X"8F5",X"8F6",X"8F7",
X"8F8",X"8F9",X"8FA",X"8FB",X"8FC",X"8FD",X"8FE",X"8FF",
X"900",X"901",X"902",X"903",X"904",X"905",X"906",X"907",
X"908",X"909",X"90A",X"90B",X"90C",X"90E",X"90F",X"910",
X"911",X"912",X"913",X"914",X"915",X"916",X"917",X"918",
X"919",X"91A",X"91C",X"91D",X"91E",X"91F",X"920",X"921",
X"922",X"923",X"924",X"925",X"926",X"928",X"929",X"92A",
X"92B",X"92C",X"92D",X"92E",X"92F",X"930",X"932",X"933",
X"934",X"935",X"936",X"937",X"938",X"93A",X"93B",X"93C",
X"93D",X"93E",X"93F",X"940",X"941",X"943",X"944",X"945",
X"946",X"947",X"948",X"94A",X"94B",X"94C",X"94D",X"94E",
X"94F",X"950",X"952",X"953",X"954",X"955",X"956",X"958",
X"959",X"95A",X"95B",X"95C",X"95D",X"95F",X"960",X"961",
X"962",X"963",X"965",X"966",X"967",X"968",X"969",X"96B",
X"96C",X"96D",X"96E",X"96F",X"971",X"972",X"973",X"974",
X"975",X"977",X"978",X"979",X"97A",X"97B",X"97D",X"97E",
X"97F",X"980",X"982",X"983",X"984",X"985",X"987",X"988",
X"989",X"98A",X"98B",X"98D",X"98E",X"98F",X"990",X"992",
X"993",X"994",X"995",X"997",X"998",X"999",X"99A",X"99C",
X"99D",X"99E",X"9A0",X"9A1",X"9A2",X"9A3",X"9A5",X"9A6",
X"9A7",X"9A8",X"9AA",X"9AB",X"9AC",X"9AE",X"9AF",X"9B0",
X"9B1",X"9B3",X"9B4",X"9B5",X"9B7",X"9B8",X"9B9",X"9BA",
X"9BC",X"9BD",X"9BE",X"9C0",X"9C1",X"9C2",X"9C3",X"9C5",
X"9C6",X"9C7",X"9C9",X"9CA",X"9CB",X"9CD",X"9CE",X"9CF",
X"9D1",X"9D2",X"9D3",X"9D5",X"9D6",X"9D7",X"9D9",X"9DA",
X"9DB",X"9DC",X"9DE",X"9DF",X"9E0",X"9E2",X"9E3",X"9E4",
X"9E6",X"9E7",X"9E8",X"9EA",X"9EB",X"9ED",X"9EE",X"9EF",
X"9F1",X"9F2",X"9F3",X"9F5",X"9F6",X"9F7",X"9F9",X"9FA",
X"9FB",X"9FD",X"9FE",X"9FF",X"A01",X"A02",X"A04",X"A05",
X"A06",X"A08",X"A09",X"A0A",X"A0C",X"A0D",X"A0E",X"A10",
X"A11",X"A13",X"A14",X"A15",X"A17",X"A18",X"A1A",X"A1B",
X"A1C",X"A1E",X"A1F",X"A20",X"A22",X"A23",X"A25",X"A26",
X"A27",X"A29",X"A2A",X"A2C",X"A2D",X"A2E",X"A30",X"A31",
X"A33",X"A34",X"A35",X"A37",X"A38",X"A3A",X"A3B",X"A3C",
X"A3E",X"A3F",X"A41",X"A42",X"A44",X"A45",X"A46",X"A48",
X"A49",X"A4B",X"A4C",X"A4D",X"A4F",X"A50",X"A52",X"A53",
X"A55",X"A56",X"A57",X"A59",X"A5A",X"A5C",X"A5D",X"A5F",
X"A60",X"A61",X"A63",X"A64",X"A66",X"A67",X"A69",X"A6A",
X"A6C",X"A6D",X"A6E",X"A70",X"A71",X"A73",X"A74",X"A76",
X"A77",X"A79",X"A7A",X"A7B",X"A7D",X"A7E",X"A80",X"A81",
X"A83",X"A84",X"A86",X"A87",X"A89",X"A8A",X"A8C",X"A8D",
X"A8E",X"A90",X"A91",X"A93",X"A94",X"A96",X"A97",X"A99",
X"A9A",X"A9C",X"A9D",X"A9F",X"AA0",X"AA2",X"AA3",X"AA5",
X"AA6",X"AA8",X"AA9",X"AAA",X"AAC",X"AAD",X"AAF",X"AB0",
X"AB2",X"AB3",X"AB5",X"AB6",X"AB8",X"AB9",X"ABB",X"ABC",
X"ABE",X"ABF",X"AC1",X"AC2",X"AC4",X"AC5",X"AC7",X"AC8",
X"ACA",X"ACB",X"ACD",X"ACE",X"AD0",X"AD1",X"AD3",X"AD4",
X"AD6",X"AD7",X"AD9",X"ADA",X"ADC",X"ADD",X"ADF",X"AE0",
X"AE2",X"AE3",X"AE5",X"AE6",X"AE8",X"AE9",X"AEB",X"AEC",
X"AEE",X"AEF",X"AF1",X"AF2",X"AF4",X"AF5",X"AF7",X"AF8",
X"AFA",X"AFC",X"AFD",X"AFF",X"B00",X"B02",X"B03",X"B05",
X"B06",X"B08",X"B09",X"B0B",X"B0C",X"B0E",X"B0F",X"B11",
X"B12",X"B14",X"B15",X"B17",X"B19",X"B1A",X"B1C",X"B1D",
X"B1F",X"B20",X"B22",X"B23",X"B25",X"B26",X"B28",X"B29",
X"B2B",X"B2C",X"B2E",X"B30",X"B31",X"B33",X"B34",X"B36",
X"B37",X"B39",X"B3A",X"B3C",X"B3D",X"B3F",X"B40",X"B42",
X"B44",X"B45",X"B47",X"B48",X"B4A",X"B4B",X"B4D",X"B4E",
X"B50",X"B51",X"B53",X"B55",X"B56",X"B58",X"B59",X"B5B",
X"B5C",X"B5E",X"B5F",X"B61",X"B63",X"B64",X"B66",X"B67",
X"B69",X"B6A",X"B6C",X"B6D",X"B6F",X"B71",X"B72",X"B74",
X"B75",X"B77",X"B78",X"B7A",X"B7B",X"B7D",X"B7F",X"B80",
X"B82",X"B83",X"B85",X"B86",X"B88",X"B89",X"B8B",X"B8D",
X"B8E",X"B90",X"B91",X"B93",X"B94",X"B96",X"B98",X"B99",
X"B9B",X"B9C",X"B9E",X"B9F",X"BA1",X"BA2",X"BA4",X"BA6",
X"BA7",X"BA9",X"BAA",X"BAC",X"BAD",X"BAF",X"BB1",X"BB2",
X"BB4",X"BB5",X"BB7",X"BB8",X"BBA",X"BBC",X"BBD",X"BBF",
X"BC0",X"BC2",X"BC3",X"BC5",X"BC6",X"BC8",X"BCA",X"BCB",
X"BCD",X"BCE",X"BD0",X"BD1",X"BD3",X"BD5",X"BD6",X"BD8",
X"BD9",X"BDB",X"BDC",X"BDE",X"BE0",X"BE1",X"BE3",X"BE4",
X"BE6",X"BE7",X"BE9",X"BEB",X"BEC",X"BEE",X"BEF",X"BF1",
X"BF2",X"BF4",X"BF6",X"BF7",X"BF9",X"BFA",X"BFC",X"BFD"
);


begin


rom_select: process (clk)
begin
  if clk'event and clk = '1' then
    if en = '1' then
   	sin_out <= SIN_ROM(conv_integer(addr));
    end if;
  end if;
end process rom_select;


end rtl;
